interface TEMP_VIF(input logic clk,input logic rst_n);

endinterface
